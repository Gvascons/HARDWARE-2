module mux4_in
	(output logic [64-1:0] f_4in,
	input logic [64-1:0] MuxA_a,MuxA_b,MuxA_c,MuxA_d,
	input logic [2:0]SelMux4);

	always_comb begin
	    	case(SelMux4) 
			0: begin
				f_4in = MuxA_a;
			end 
	
			1: begin
				f_4in = MuxA_b;
			end
	
			2: begin
				f_4in = MuxA_c;
			end 
			3: begin
				f_4in = MuxA_d;
			end 
		endcase 
	end
endmodule